module sample_test ();
    initial begin
        $display(3 == 3);
    end
endmodule