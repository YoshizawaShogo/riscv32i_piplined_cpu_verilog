module hello_test;

    initial begin
        $display("Hello world 2");
    end
endmodule