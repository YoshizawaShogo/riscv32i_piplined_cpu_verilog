module hello_test;

    initial begin
        $display("Hello world");
    end
endmodule