// RV32Iのみ(例外処理もなし)

// alu fn
`define ALU_FN_LEN 4
`define ALU_X    `ALU_FN_LEN'd0
`define ALU_ADD  `ALU_FN_LEN'd1
`define ALU_SUB  `ALU_FN_LEN'd2
`define ALU_AND  `ALU_FN_LEN'd3
`define ALU_OR   `ALU_FN_LEN'd4
`define ALU_XOR  `ALU_FN_LEN'd5
`define ALU_SLL  `ALU_FN_LEN'd6
`define ALU_SRL  `ALU_FN_LEN'd7
`define ALU_SRA  `ALU_FN_LEN'd8
`define ALU_SLT  `ALU_FN_LEN'd9
`define ALU_SLTU `ALU_FN_LEN'd10
`define ALU_JALR `ALU_FN_LEN'd11

// branch fn
`define BR_FN_LEN 3
`define BR_X     `BR_FN_LEN'd0
`define BR_BEQ   `BR_FN_LEN'd1
`define BR_BNE   `BR_FN_LEN'd2
`define BR_BLT   `BR_FN_LEN'd3
`define BR_BGE   `BR_FN_LEN'd4
`define BR_BLTU  `BR_FN_LEN'd5
`define BR_BGEU  `BR_FN_LEN'd6
`define BR_JAL   `BR_FN_LEN'd7

// rs1
`define RS1_LEN 2
`define RS1_X    `RS1_LEN'd0
`define RS1_RS1  `RS1_LEN'd1
`define RS1_PC   `RS1_LEN'd2

// rs2
`define RS2_LEN 2
`define RS2_X    `RS2_LEN'd0
`define RS2_RS2  `RS2_LEN'd1
`define RS2_IMI  `RS2_LEN'd2

// mem_fn
`define MEM_FN_LEN 3
`define MEM_LB   `MEM_FN_LEN'd0
`define MEM_LH   `MEM_FN_LEN'd1
`define MEM_LW   `MEM_FN_LEN'd2
`define MEM_LBU  `MEM_FN_LEN'd3
`define MEM_LHU  `MEM_FN_LEN'd4
`define MEM_SB   `MEM_FN_LEN'd5
`define MEM_SH   `MEM_FN_LEN'd6
`define MEM_SW   `MEM_FN_LEN'd7

// wb_sel
`define WB_FN_LEN 2
`define WB_X      `WB_FN_LEN'd0
`define WB_ALU    `WB_FN_LEN'd1
`define WB_MEM    `WB_FN_LEN'd2
`define WB_PC     `WB_FN_LEN'd3

// ecall
`define ECALL_FLAG_LEN 1
`define ECALL_N `ECALL_FLAG_LEN'b0
`define ECALL_Y `ECALL_FLAG_LEN'b1

/* 以下命令コード */
// https://riscv.org/wp-content/uploads/2017/05/riscv-spec-v2.2.pdf の p.116参照
// ロード・ストア
`define LUI     32'b?????????????????????????0110111
`define AUIPC   32'b?????????????????????????0010111
`define JAL     32'b?????????????????????????1101111
`define JALR    32'b?????????????????000?????1100111
`define BEQ     32'b?????????????????000?????1100011
`define BNE     32'b?????????????????001?????1100011
`define BLT     32'b?????????????????100?????1100011
`define BGE     32'b?????????????????101?????1100011
`define BLTU    32'b?????????????????110?????1100011
`define BGEU    32'b?????????????????111?????1100011
`define LB      32'b?????????????????000?????0000011
`define LH      32'b?????????????????001?????0000011
`define LW      32'b?????????????????010?????0000011
`define LBU     32'b?????????????????100?????0000011
`define LHU     32'b?????????????????101?????0000011
`define SB      32'b?????????????????000?????0100011
`define SH      32'b?????????????????001?????0100011
`define SW      32'b?????????????????010?????0100011
`define ADDI    32'b?????????????????000?????0010011
`define SLTI    32'b?????????????????010?????0010011
`define SLTIU   32'b?????????????????011?????0010011
`define XORI    32'b?????????????????100?????0010011
`define ORI     32'b?????????????????110?????0010011
`define ANDI    32'b?????????????????111?????0010011
`define SLLI    32'b0000000??????????001?????0010011
`define SRLI    32'b0000000??????????101?????0010011
`define SRAI    32'b0100000??????????101?????0010011
`define ADD     32'b0000000??????????000?????0110011
`define SUB     32'b0100000??????????000?????0110011
`define SLL     32'b0000000??????????001?????0110011
`define SLT     32'b0000000??????????010?????0110011
`define SLTU    32'b0000000??????????011?????0110011
`define XOR     32'b0000000??????????100?????0110011
`define SRL     32'b0000000??????????101?????0110011
`define SRA     32'b0100000??????????101?????0110011
`define OR      32'b0000000??????????110?????0110011
`define AND     32'b0000000??????????111?????0110011
`define FENCE   32'b0000????????00000000000000001111
`define FENCE_I 32'b00000000000000000001000000001111
`define ECALL   32'b00000000000000000000000001110011
`define CSRRW   32'??????????????????001?????1110011
`define CSRRS   32'??????????????????010?????1110011
`define CSRRC   32'??????????????????011?????1110011
`define CSRRWI  32'??????????????????101?????1110011
`define CSRRSI  32'??????????????????110?????1110011
`define CSRRCI  32'??????????????????111?????1110011